module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _112_;
 wire _113_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire \dpath/a_lt_b$in0[10] ;
 wire \dpath/a_lt_b$in0[11] ;
 wire \dpath/a_lt_b$in0[12] ;
 wire \dpath/a_lt_b$in0[13] ;
 wire \dpath/a_lt_b$in0[14] ;
 wire \dpath/a_lt_b$in0[15] ;
 wire \dpath/a_lt_b$in0[1] ;
 wire \dpath/a_lt_b$in0[2] ;
 wire \dpath/a_lt_b$in0[3] ;
 wire \dpath/a_lt_b$in0[4] ;
 wire \dpath/a_lt_b$in0[5] ;
 wire \dpath/a_lt_b$in0[6] ;
 wire \dpath/a_lt_b$in0[7] ;
 wire \dpath/a_lt_b$in0[8] ;
 wire \dpath/a_lt_b$in0[9] ;
 wire \dpath/a_lt_b$in1[0] ;
 wire \dpath/a_lt_b$in1[1] ;
 wire cut_1911;
 wire cut_1922;
 wire cut_1933;
 wire cut_1944;
 wire cut_1955;
 wire cut_1966;
 wire cut_1977;
 wire cut_1988;
 wire cut_1999;
 wire cut_20010;
 wire cut_20111;
 wire cut_20212;
 wire cut_20313;
 wire cut_20414;
 wire cut_20515;
 wire cut_20616;
 wire cut_20717;
 wire cut_20818;
 wire cut_20919;
 wire cut_21020;
 wire cut_21121;
 wire cut_21222;
 wire cut_21323;
 wire cut_21424;
 wire cut_21525;
 wire cut_21626;
 wire cut_21727;
 wire cut_21828;
 wire cut_21929;
 wire cut_22030;
 wire cut_22131;
 wire cut_22232;
 wire cut_22333;
 wire cut_22434;
 wire cut_22535;
 wire cut_22636;
 wire cut_22737;
 wire cut_22838;
 wire cut_22939;
 wire cut_23040;
 wire cut_23141;
 wire cut_23242;
 wire cut_23343;
 wire cut_23444;
 wire cut_23545;
 wire cut_23646;
 wire cut_23747;
 wire cut_23848;
 wire cut_23949;
 wire cut_24050;
 wire cut_24151;
 wire cut_24252;
 wire cut_24353;
 wire cut_24454;
 wire cut_24555;
 wire cut_24656;
 wire cut_24757;
 wire cut_24858;
 wire cut_24959;
 wire cut_25060;
 wire cut_25161;
 wire cut_25262;
 wire cut_25363;
 wire cut_25464;
 wire cut_25565;
 wire cut_25666;
 wire cut_25767;
 wire cut_25868;
 wire cut_25969;
 wire cut_26070;
 wire cut_26171;
 wire cut_26272;
 wire cut_26373;
 wire cut_26474;
 wire cut_26575;
 wire cut_26676;
 wire cut_26777;
 wire cut_26878;
 wire cut_26979;
 wire cut_27080;
 wire cut_27181;
 wire cut_27282;
 wire cut_27383;
 wire cut_27484;
 wire cut_27585;
 wire cut_27686;
 wire cut_27787;
 wire cut_27888;
 wire cut_27989;
 wire cut_28090;
 wire cut_28191;
 wire cut_28292;
 wire cut_28393;
 wire cut_28494;
 wire cut_28595;
 wire cut_28696;
 wire cut_28797;
 wire cut_28898;
 wire cut_28999;
 wire cut_290100;
 wire cut_291101;
 wire cut_292102;
 wire cut_293103;
 wire cut_294104;
 wire cut_295105;
 wire cut_296106;
 wire cut_297107;
 wire cut_298108;
 wire cut_299109;
 wire cut_300110;
 wire cut_301111;
 wire cut_302112;
 wire cut_303113;
 wire cut_304114;
 wire cut_305115;
 wire cut_306116;
 wire cut_307117;
 wire cut_308118;
 wire cut_309119;
 wire cut_310120;
 wire cut_311121;

 INVx1_ASAP7_75t_R _259_ (.A(req_val),
    .Y(_112_));
 AO21x1_ASAP7_75t_R _261_ (.A1(_112_),
    .A2(req_rdy),
    .B(_113_),
    .Y(_000_));
 FAx1_ASAP7_75t_R _420_ (.SN(_030_),
    .A(_208_),
    .B(\dpath/a_lt_b$in1[1] ),
    .CI(_209_),
    .CON(_028_));
 HAxp5_ASAP7_75t_R _421_ (.A(\dpath/a_lt_b$in1[0] ),
    .B(_210_),
    .CON(_226_),
    .SN(resp_msg[0]));
 HAxp5_ASAP7_75t_R _422_ (.A(_211_),
    .B(\dpath/a_lt_b$in0[15] ),
    .CON(_003_),
    .SN(_048_));
 HAxp5_ASAP7_75t_R _423_ (.A(_212_),
    .B(\dpath/a_lt_b$in0[14] ),
    .CON(_004_),
    .SN(_005_));
 HAxp5_ASAP7_75t_R _424_ (.A(_213_),
    .B(\dpath/a_lt_b$in0[13] ),
    .CON(_006_),
    .SN(_007_));
 HAxp5_ASAP7_75t_R _425_ (.A(_214_),
    .B(\dpath/a_lt_b$in0[12] ),
    .CON(_008_),
    .SN(_009_));
 HAxp5_ASAP7_75t_R _426_ (.A(_215_),
    .B(\dpath/a_lt_b$in0[11] ),
    .CON(_010_),
    .SN(_011_));
 HAxp5_ASAP7_75t_R _427_ (.A(_216_),
    .B(\dpath/a_lt_b$in0[10] ),
    .CON(_012_),
    .SN(_013_));
 HAxp5_ASAP7_75t_R _428_ (.A(_217_),
    .B(\dpath/a_lt_b$in0[9] ),
    .CON(_014_),
    .SN(_049_));
 HAxp5_ASAP7_75t_R _429_ (.A(_218_),
    .B(\dpath/a_lt_b$in0[8] ),
    .CON(_015_),
    .SN(_016_));
 HAxp5_ASAP7_75t_R _430_ (.A(_219_),
    .B(\dpath/a_lt_b$in0[7] ),
    .CON(_017_),
    .SN(_050_));
 HAxp5_ASAP7_75t_R _431_ (.A(_220_),
    .B(\dpath/a_lt_b$in0[6] ),
    .CON(_018_),
    .SN(_019_));
 HAxp5_ASAP7_75t_R _432_ (.A(_221_),
    .B(\dpath/a_lt_b$in0[5] ),
    .CON(_020_),
    .SN(_051_));
 HAxp5_ASAP7_75t_R _433_ (.A(_222_),
    .B(\dpath/a_lt_b$in0[4] ),
    .CON(_021_),
    .SN(_022_));
 HAxp5_ASAP7_75t_R _434_ (.A(_223_),
    .B(\dpath/a_lt_b$in0[3] ),
    .CON(_023_),
    .SN(_024_));
 HAxp5_ASAP7_75t_R _435_ (.A(_224_),
    .B(\dpath/a_lt_b$in0[2] ),
    .CON(_025_),
    .SN(_026_));
 HAxp5_ASAP7_75t_R _436_ (.A(_225_),
    .B(\dpath/a_lt_b$in0[1] ),
    .CON(_027_),
    .SN(_052_));
 DFFHQNx1_ASAP7_75t_R \ctrl/state/out[1]$_DFF_P_  (.CLK(clk),
    .D(_001_),
    .QN(_047_));
 DFFHQNx1_ASAP7_75t_R \ctrl/state/out[2]$_DFF_P_  (.CLK(clk),
    .D(_002_),
    .QN(_046_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[0]$_DFFE_PP_  (.CLK(clk),
    .D(_069_),
    .QN(_210_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[10]$_DFFE_PP_  (.CLK(clk),
    .D(_079_),
    .QN(_036_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[11]$_DFFE_PP_  (.CLK(clk),
    .D(_080_),
    .QN(_035_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[12]$_DFFE_PP_  (.CLK(clk),
    .D(_081_),
    .QN(_034_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[13]$_DFFE_PP_  (.CLK(clk),
    .D(_082_),
    .QN(_033_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[14]$_DFFE_PP_  (.CLK(clk),
    .D(_083_),
    .QN(_032_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[15]$_DFFE_PP_  (.CLK(clk),
    .D(_084_),
    .QN(_031_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[1]$_DFFE_PP_  (.CLK(clk),
    .D(_070_),
    .QN(_209_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[2]$_DFFE_PP_  (.CLK(clk),
    .D(_071_),
    .QN(_044_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[3]$_DFFE_PP_  (.CLK(clk),
    .D(_072_),
    .QN(_043_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[4]$_DFFE_PP_  (.CLK(clk),
    .D(_073_),
    .QN(_042_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[5]$_DFFE_PP_  (.CLK(clk),
    .D(_074_),
    .QN(_041_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[6]$_DFFE_PP_  (.CLK(clk),
    .D(_075_),
    .QN(_040_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[7]$_DFFE_PP_  (.CLK(clk),
    .D(_076_),
    .QN(_039_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[8]$_DFFE_PP_  (.CLK(clk),
    .D(_077_),
    .QN(_038_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in0[9]$_DFFE_PP_  (.CLK(clk),
    .D(_078_),
    .QN(_037_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[0]$_DFFE_PP_  (.CLK(clk),
    .D(_053_),
    .QN(_045_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[10]$_DFFE_PP_  (.CLK(clk),
    .D(_063_),
    .QN(_216_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[11]$_DFFE_PP_  (.CLK(clk),
    .D(_064_),
    .QN(_215_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[12]$_DFFE_PP_  (.CLK(clk),
    .D(_065_),
    .QN(_214_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[13]$_DFFE_PP_  (.CLK(clk),
    .D(_066_),
    .QN(_213_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[14]$_DFFE_PP_  (.CLK(clk),
    .D(_067_),
    .QN(_212_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[15]$_DFFE_PP_  (.CLK(clk),
    .D(_068_),
    .QN(_211_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[1]$_DFFE_PP_  (.CLK(clk),
    .D(_054_),
    .QN(_225_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[2]$_DFFE_PP_  (.CLK(clk),
    .D(_055_),
    .QN(_224_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[3]$_DFFE_PP_  (.CLK(clk),
    .D(_056_),
    .QN(_223_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[4]$_DFFE_PP_  (.CLK(clk),
    .D(_057_),
    .QN(_222_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[5]$_DFFE_PP_  (.CLK(clk),
    .D(_058_),
    .QN(_221_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[6]$_DFFE_PP_  (.CLK(clk),
    .D(_059_),
    .QN(_220_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[7]$_DFFE_PP_  (.CLK(clk),
    .D(_060_),
    .QN(_219_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[8]$_DFFE_PP_  (.CLK(clk),
    .D(_061_),
    .QN(_218_));
 DFFHQNx1_ASAP7_75t_R \dpath/a_lt_b$in1[9]$_DFFE_PP_  (.CLK(clk),
    .D(_062_),
    .QN(_217_));
 DFFHQNx1_ASAP7_75t_R \req_rdy$_DFF_P_  (.CLK(clk),
    .D(_000_),
    .QN(_029_));
 INVx1_ASAP7_75t_R cut_0 (.A(_225_),
    .Y(\dpath/a_lt_b$in1[1] ));
 INVx1_ASAP7_75t_R cut_1 (.A(_045_),
    .Y(\dpath/a_lt_b$in1[0] ));
 BUFx2_ASAP7_75t_R cut_2 (.A(_029_),
    .Y(cut_1911));
 INVx1_ASAP7_75t_R cut_3 (.A(cut_1911),
    .Y(cut_1922));
 BUFx2_ASAP7_75t_R cut_4 (.A(cut_1922),
    .Y(req_rdy));
 INVx1_ASAP7_75t_R cut_5 (.A(reset),
    .Y(cut_21424));
 NOR2x1_ASAP7_75t_R cut_6 (.A(reset),
    .B(_046_),
    .Y(cut_21525));
 INVx1_ASAP7_75t_R cut_7 (.A(_028_),
    .Y(cut_1933));
 OA21x2_ASAP7_75t_R cut_8 (.A1(_026_),
    .A2(cut_1933),
    .B(_025_),
    .Y(cut_1944));
 OA21x2_ASAP7_75t_R cut_9 (.A1(_024_),
    .A2(cut_1944),
    .B(_023_),
    .Y(cut_1955));
 OA21x2_ASAP7_75t_R cut_10 (.A1(_022_),
    .A2(cut_1955),
    .B(_021_),
    .Y(cut_1966));
 OA21x2_ASAP7_75t_R cut_11 (.A1(_051_),
    .A2(cut_1966),
    .B(_020_),
    .Y(cut_1977));
 OA21x2_ASAP7_75t_R cut_12 (.A1(_019_),
    .A2(cut_1977),
    .B(_018_),
    .Y(cut_1988));
 OA21x2_ASAP7_75t_R cut_13 (.A1(_050_),
    .A2(cut_1988),
    .B(_017_),
    .Y(cut_1999));
 OA21x2_ASAP7_75t_R cut_14 (.A1(_016_),
    .A2(cut_1999),
    .B(_015_),
    .Y(cut_20010));
 OA21x2_ASAP7_75t_R cut_15 (.A1(_049_),
    .A2(cut_20010),
    .B(_014_),
    .Y(cut_20111));
 OA21x2_ASAP7_75t_R cut_16 (.A1(_013_),
    .A2(cut_20111),
    .B(_012_),
    .Y(cut_20212));
 OA21x2_ASAP7_75t_R cut_17 (.A1(_011_),
    .A2(cut_20212),
    .B(_010_),
    .Y(cut_20313));
 OA21x2_ASAP7_75t_R cut_18 (.A1(_009_),
    .A2(cut_20313),
    .B(_008_),
    .Y(cut_20414));
 OA21x2_ASAP7_75t_R cut_19 (.A1(_007_),
    .A2(cut_20414),
    .B(_006_),
    .Y(cut_20515));
 OA21x2_ASAP7_75t_R cut_20 (.A1(_005_),
    .A2(cut_20515),
    .B(_004_),
    .Y(cut_20616));
 OAI21x1_ASAP7_75t_R cut_21 (.A1(_048_),
    .A2(cut_20616),
    .B(_003_),
    .Y(cut_20717));
 BUFx2_ASAP7_75t_R cut_22 (.A(cut_20717),
    .Y(cut_21222));
 AND4x1_ASAP7_75t_R cut_23 (.A(_215_),
    .B(_216_),
    .C(_217_),
    .D(_218_),
    .Y(cut_20818));
 AND4x1_ASAP7_75t_R cut_24 (.A(_211_),
    .B(_212_),
    .C(_213_),
    .D(_214_),
    .Y(cut_20919));
 AND4x1_ASAP7_75t_R cut_25 (.A(_223_),
    .B(_224_),
    .C(_225_),
    .D(_045_),
    .Y(cut_21020));
 AND4x1_ASAP7_75t_R cut_26 (.A(_219_),
    .B(_220_),
    .C(_221_),
    .D(_222_),
    .Y(cut_21121));
 AND4x1_ASAP7_75t_R cut_27 (.A(cut_20818),
    .B(cut_20919),
    .C(cut_21020),
    .D(cut_21121),
    .Y(cut_21323));
 NAND2x1_ASAP7_75t_R cut_28 (.A(cut_21222),
    .B(cut_21323),
    .Y(cut_21626));
 AO32x1_ASAP7_75t_R cut_29 (.A1(cut_21424),
    .A2(req_val),
    .A3(req_rdy),
    .B1(cut_21525),
    .B2(cut_21626),
    .Y(_002_));
 INVx1_ASAP7_75t_R cut_30 (.A(_047_),
    .Y(cut_21727));
 AND3x1_ASAP7_75t_R cut_31 (.A(cut_1911),
    .B(_046_),
    .C(cut_21727),
    .Y(resp_val));
 AO21x1_ASAP7_75t_R cut_32 (.A1(resp_rdy),
    .A2(resp_val),
    .B(reset),
    .Y(_113_));
 OR2x2_ASAP7_75t_R cut_33 (.A(reset),
    .B(_046_),
    .Y(cut_21828));
 OAI22x1_ASAP7_75t_R cut_34 (.A1(cut_21828),
    .A2(cut_21626),
    .B1(_113_),
    .B2(_047_),
    .Y(_001_));
 INVx1_ASAP7_75t_R cut_35 (.A(_031_),
    .Y(\dpath/a_lt_b$in0[15] ));
 INVx1_ASAP7_75t_R cut_36 (.A(_032_),
    .Y(\dpath/a_lt_b$in0[14] ));
 INVx1_ASAP7_75t_R cut_37 (.A(_033_),
    .Y(\dpath/a_lt_b$in0[13] ));
 INVx1_ASAP7_75t_R cut_38 (.A(_034_),
    .Y(\dpath/a_lt_b$in0[12] ));
 INVx1_ASAP7_75t_R cut_39 (.A(_035_),
    .Y(\dpath/a_lt_b$in0[11] ));
 INVx1_ASAP7_75t_R cut_40 (.A(_036_),
    .Y(\dpath/a_lt_b$in0[10] ));
 INVx1_ASAP7_75t_R cut_41 (.A(_037_),
    .Y(\dpath/a_lt_b$in0[9] ));
 INVx1_ASAP7_75t_R cut_42 (.A(_038_),
    .Y(\dpath/a_lt_b$in0[8] ));
 INVx1_ASAP7_75t_R cut_43 (.A(_039_),
    .Y(\dpath/a_lt_b$in0[7] ));
 INVx1_ASAP7_75t_R cut_44 (.A(_040_),
    .Y(\dpath/a_lt_b$in0[6] ));
 INVx1_ASAP7_75t_R cut_45 (.A(_041_),
    .Y(\dpath/a_lt_b$in0[5] ));
 INVx1_ASAP7_75t_R cut_46 (.A(_042_),
    .Y(\dpath/a_lt_b$in0[4] ));
 INVx1_ASAP7_75t_R cut_47 (.A(_043_),
    .Y(\dpath/a_lt_b$in0[3] ));
 INVx1_ASAP7_75t_R cut_48 (.A(_044_),
    .Y(\dpath/a_lt_b$in0[2] ));
 INVx1_ASAP7_75t_R cut_49 (.A(_209_),
    .Y(\dpath/a_lt_b$in0[1] ));
 BUFx2_ASAP7_75t_R cut_50 (.A(cut_1922),
    .Y(cut_22333));
 OA21x2_ASAP7_75t_R cut_51 (.A1(_046_),
    .A2(cut_20717),
    .B(cut_1911),
    .Y(cut_21929));
 BUFx2_ASAP7_75t_R cut_52 (.A(cut_21929),
    .Y(cut_22434));
 INVx1_ASAP7_75t_R cut_53 (.A(_046_),
    .Y(cut_22030));
 AND2x2_ASAP7_75t_R cut_54 (.A(_029_),
    .B(cut_22030),
    .Y(cut_22131));
 OA211x2_ASAP7_75t_R cut_55 (.A1(_048_),
    .A2(cut_20616),
    .B(cut_22131),
    .C(_003_),
    .Y(cut_22232));
 BUFx2_ASAP7_75t_R cut_56 (.A(cut_22232),
    .Y(cut_22535));
 INVx1_ASAP7_75t_R cut_57 (.A(_210_),
    .Y(cut_22636));
 AO222x2_ASAP7_75t_R cut_58 (.A1(cut_22333),
    .A2(req_msg[0]),
    .B1(cut_22434),
    .B2(\dpath/a_lt_b$in1[0] ),
    .C1(cut_22535),
    .C2(cut_22636),
    .Y(_053_));
 BUFx2_ASAP7_75t_R cut_59 (.A(cut_1922),
    .Y(cut_22737));
 AO222x2_ASAP7_75t_R cut_60 (.A1(cut_22737),
    .A2(req_msg[1]),
    .B1(cut_22434),
    .B2(\dpath/a_lt_b$in1[1] ),
    .C1(cut_22535),
    .C2(\dpath/a_lt_b$in0[1] ),
    .Y(_054_));
 INVx1_ASAP7_75t_R cut_61 (.A(_224_),
    .Y(cut_22838));
 AO222x2_ASAP7_75t_R cut_62 (.A1(cut_22737),
    .A2(req_msg[2]),
    .B1(cut_22434),
    .B2(cut_22838),
    .C1(cut_22535),
    .C2(\dpath/a_lt_b$in0[2] ),
    .Y(_055_));
 INVx1_ASAP7_75t_R cut_63 (.A(_223_),
    .Y(cut_22939));
 AO222x2_ASAP7_75t_R cut_64 (.A1(cut_22737),
    .A2(req_msg[3]),
    .B1(cut_22434),
    .B2(cut_22939),
    .C1(cut_22535),
    .C2(\dpath/a_lt_b$in0[3] ),
    .Y(_056_));
 INVx1_ASAP7_75t_R cut_65 (.A(_222_),
    .Y(cut_23040));
 AO222x2_ASAP7_75t_R cut_66 (.A1(cut_22737),
    .A2(req_msg[4]),
    .B1(cut_22434),
    .B2(cut_23040),
    .C1(cut_22535),
    .C2(\dpath/a_lt_b$in0[4] ),
    .Y(_057_));
 INVx1_ASAP7_75t_R cut_67 (.A(_221_),
    .Y(cut_23141));
 AO222x2_ASAP7_75t_R cut_68 (.A1(cut_22737),
    .A2(req_msg[5]),
    .B1(cut_22434),
    .B2(cut_23141),
    .C1(cut_22535),
    .C2(\dpath/a_lt_b$in0[5] ),
    .Y(_058_));
 INVx1_ASAP7_75t_R cut_69 (.A(_220_),
    .Y(cut_23242));
 AO222x2_ASAP7_75t_R cut_70 (.A1(cut_22737),
    .A2(req_msg[6]),
    .B1(cut_22434),
    .B2(cut_23242),
    .C1(cut_22535),
    .C2(\dpath/a_lt_b$in0[6] ),
    .Y(_059_));
 INVx1_ASAP7_75t_R cut_71 (.A(_219_),
    .Y(cut_23343));
 AO222x2_ASAP7_75t_R cut_72 (.A1(cut_22737),
    .A2(req_msg[7]),
    .B1(cut_22434),
    .B2(cut_23343),
    .C1(cut_22535),
    .C2(\dpath/a_lt_b$in0[7] ),
    .Y(_060_));
 INVx1_ASAP7_75t_R cut_73 (.A(_218_),
    .Y(cut_23444));
 AO222x2_ASAP7_75t_R cut_74 (.A1(cut_22737),
    .A2(req_msg[8]),
    .B1(cut_22434),
    .B2(cut_23444),
    .C1(cut_22535),
    .C2(\dpath/a_lt_b$in0[8] ),
    .Y(_061_));
 INVx1_ASAP7_75t_R cut_75 (.A(_217_),
    .Y(cut_23545));
 AO222x2_ASAP7_75t_R cut_76 (.A1(cut_22737),
    .A2(req_msg[9]),
    .B1(cut_22434),
    .B2(cut_23545),
    .C1(cut_22535),
    .C2(\dpath/a_lt_b$in0[9] ),
    .Y(_062_));
 INVx1_ASAP7_75t_R cut_77 (.A(_216_),
    .Y(cut_23646));
 BUFx2_ASAP7_75t_R cut_78 (.A(cut_22232),
    .Y(cut_23747));
 AO222x2_ASAP7_75t_R cut_79 (.A1(cut_22737),
    .A2(req_msg[10]),
    .B1(cut_21929),
    .B2(cut_23646),
    .C1(cut_23747),
    .C2(\dpath/a_lt_b$in0[10] ),
    .Y(_063_));
 INVx1_ASAP7_75t_R cut_80 (.A(_215_),
    .Y(cut_23848));
 AO222x2_ASAP7_75t_R cut_81 (.A1(cut_1922),
    .A2(req_msg[11]),
    .B1(cut_21929),
    .B2(cut_23848),
    .C1(cut_23747),
    .C2(\dpath/a_lt_b$in0[11] ),
    .Y(_064_));
 INVx1_ASAP7_75t_R cut_82 (.A(_214_),
    .Y(cut_23949));
 AO222x2_ASAP7_75t_R cut_83 (.A1(cut_1922),
    .A2(req_msg[12]),
    .B1(cut_21929),
    .B2(cut_23949),
    .C1(cut_23747),
    .C2(\dpath/a_lt_b$in0[12] ),
    .Y(_065_));
 INVx1_ASAP7_75t_R cut_84 (.A(_213_),
    .Y(cut_24050));
 AO222x2_ASAP7_75t_R cut_85 (.A1(cut_1922),
    .A2(req_msg[13]),
    .B1(cut_21929),
    .B2(cut_24050),
    .C1(cut_23747),
    .C2(\dpath/a_lt_b$in0[13] ),
    .Y(_066_));
 INVx1_ASAP7_75t_R cut_86 (.A(_212_),
    .Y(cut_24151));
 AO222x2_ASAP7_75t_R cut_87 (.A1(cut_1922),
    .A2(req_msg[14]),
    .B1(cut_21929),
    .B2(cut_24151),
    .C1(cut_23747),
    .C2(\dpath/a_lt_b$in0[14] ),
    .Y(_067_));
 INVx1_ASAP7_75t_R cut_88 (.A(_211_),
    .Y(cut_24252));
 AO222x2_ASAP7_75t_R cut_89 (.A1(cut_1922),
    .A2(req_msg[15]),
    .B1(cut_21929),
    .B2(cut_24252),
    .C1(cut_23747),
    .C2(\dpath/a_lt_b$in0[15] ),
    .Y(_068_));
 BUFx2_ASAP7_75t_R cut_90 (.A(cut_22030),
    .Y(cut_24656));
 AND3x1_ASAP7_75t_R cut_91 (.A(resp_msg[0]),
    .B(cut_20717),
    .C(cut_22131),
    .Y(cut_24757));
 BUFx2_ASAP7_75t_R cut_92 (.A(cut_1911),
    .Y(cut_24454));
 NAND2x1_ASAP7_75t_R cut_93 (.A(_029_),
    .B(cut_22030),
    .Y(cut_24353));
 BUFx2_ASAP7_75t_R cut_94 (.A(cut_24353),
    .Y(cut_24555));
 OA21x2_ASAP7_75t_R cut_95 (.A1(cut_24454),
    .A2(req_msg[16]),
    .B(cut_24555),
    .Y(cut_24858));
 AND2x2_ASAP7_75t_R cut_96 (.A(\dpath/a_lt_b$in1[0] ),
    .B(cut_23747),
    .Y(cut_24959));
 OA33x2_ASAP7_75t_R cut_97 (.A1(req_rdy),
    .A2(cut_22636),
    .A3(cut_24656),
    .B1(cut_24757),
    .B2(cut_24858),
    .B3(cut_24959),
    .Y(_069_));
 INVx1_ASAP7_75t_R cut_98 (.A(_030_),
    .Y(resp_msg[1]));
 AND3x1_ASAP7_75t_R cut_99 (.A(resp_msg[1]),
    .B(cut_20717),
    .C(cut_22131),
    .Y(cut_25060));
 OA21x2_ASAP7_75t_R cut_100 (.A1(cut_24454),
    .A2(req_msg[17]),
    .B(cut_24555),
    .Y(cut_25161));
 AND2x2_ASAP7_75t_R cut_101 (.A(\dpath/a_lt_b$in1[1] ),
    .B(cut_23747),
    .Y(cut_25262));
 OA33x2_ASAP7_75t_R cut_102 (.A1(req_rdy),
    .A2(\dpath/a_lt_b$in0[1] ),
    .A3(cut_24656),
    .B1(cut_25060),
    .B2(cut_25161),
    .B3(cut_25262),
    .Y(_070_));
 BUFx2_ASAP7_75t_R cut_103 (.A(cut_22232),
    .Y(cut_25363));
 AND2x2_ASAP7_75t_R cut_104 (.A(cut_22838),
    .B(cut_25363),
    .Y(cut_25565));
 OA21x2_ASAP7_75t_R cut_105 (.A1(cut_24454),
    .A2(req_msg[18]),
    .B(cut_24555),
    .Y(cut_25666));
 BUFx2_ASAP7_75t_R cut_106 (.A(cut_22131),
    .Y(cut_25464));
 XNOR2x2_ASAP7_75t_R cut_107 (.A(_026_),
    .B(_028_),
    .Y(resp_msg[2]));
 AND3x1_ASAP7_75t_R cut_108 (.A(cut_21222),
    .B(cut_25464),
    .C(resp_msg[2]),
    .Y(cut_25767));
 OA33x2_ASAP7_75t_R cut_109 (.A1(req_rdy),
    .A2(\dpath/a_lt_b$in0[2] ),
    .A3(cut_24656),
    .B1(cut_25565),
    .B2(cut_25666),
    .B3(cut_25767),
    .Y(_071_));
 AND2x2_ASAP7_75t_R cut_110 (.A(cut_22939),
    .B(cut_25363),
    .Y(cut_26070));
 OA21x2_ASAP7_75t_R cut_111 (.A1(cut_24454),
    .A2(req_msg[19]),
    .B(cut_24555),
    .Y(cut_26171));
 INVx1_ASAP7_75t_R cut_112 (.A(_226_),
    .Y(_208_));
 OA21x2_ASAP7_75t_R cut_113 (.A1(_208_),
    .A2(_052_),
    .B(_027_),
    .Y(cut_25868));
 OA21x2_ASAP7_75t_R cut_114 (.A1(_026_),
    .A2(cut_25868),
    .B(_025_),
    .Y(cut_25969));
 XOR2x2_ASAP7_75t_R cut_115 (.A(_024_),
    .B(cut_25969),
    .Y(resp_msg[3]));
 AND3x1_ASAP7_75t_R cut_116 (.A(cut_21222),
    .B(cut_25464),
    .C(resp_msg[3]),
    .Y(cut_26272));
 OA33x2_ASAP7_75t_R cut_117 (.A1(req_rdy),
    .A2(\dpath/a_lt_b$in0[3] ),
    .A3(cut_24656),
    .B1(cut_26070),
    .B2(cut_26171),
    .B3(cut_26272),
    .Y(_072_));
 XOR2x2_ASAP7_75t_R cut_118 (.A(_022_),
    .B(cut_1955),
    .Y(resp_msg[4]));
 AND3x1_ASAP7_75t_R cut_119 (.A(cut_20717),
    .B(cut_22131),
    .C(resp_msg[4]),
    .Y(cut_26373));
 OA21x2_ASAP7_75t_R cut_120 (.A1(cut_24454),
    .A2(req_msg[20]),
    .B(cut_24555),
    .Y(cut_26474));
 AND2x2_ASAP7_75t_R cut_121 (.A(cut_23040),
    .B(cut_23747),
    .Y(cut_26575));
 OA33x2_ASAP7_75t_R cut_122 (.A1(req_rdy),
    .A2(\dpath/a_lt_b$in0[4] ),
    .A3(cut_24656),
    .B1(cut_26373),
    .B2(cut_26474),
    .B3(cut_26575),
    .Y(_073_));
 AND2x2_ASAP7_75t_R cut_123 (.A(cut_23141),
    .B(cut_25363),
    .Y(cut_26878));
 OA21x2_ASAP7_75t_R cut_124 (.A1(cut_24454),
    .A2(req_msg[21]),
    .B(cut_24555),
    .Y(cut_26979));
 OA21x2_ASAP7_75t_R cut_125 (.A1(_024_),
    .A2(cut_25969),
    .B(_023_),
    .Y(cut_26676));
 OA21x2_ASAP7_75t_R cut_126 (.A1(_022_),
    .A2(cut_26676),
    .B(_021_),
    .Y(cut_26777));
 XOR2x2_ASAP7_75t_R cut_127 (.A(_051_),
    .B(cut_26777),
    .Y(resp_msg[5]));
 AND3x1_ASAP7_75t_R cut_128 (.A(cut_21222),
    .B(cut_25464),
    .C(resp_msg[5]),
    .Y(cut_27080));
 OA33x2_ASAP7_75t_R cut_129 (.A1(req_rdy),
    .A2(\dpath/a_lt_b$in0[5] ),
    .A3(cut_24656),
    .B1(cut_26878),
    .B2(cut_26979),
    .B3(cut_27080),
    .Y(_074_));
 AND2x2_ASAP7_75t_R cut_130 (.A(cut_23242),
    .B(cut_25363),
    .Y(cut_27181));
 OA21x2_ASAP7_75t_R cut_131 (.A1(cut_24454),
    .A2(req_msg[22]),
    .B(cut_24555),
    .Y(cut_27282));
 XOR2x2_ASAP7_75t_R cut_132 (.A(_019_),
    .B(cut_1977),
    .Y(resp_msg[6]));
 AND3x1_ASAP7_75t_R cut_133 (.A(cut_21222),
    .B(cut_25464),
    .C(resp_msg[6]),
    .Y(cut_27383));
 OA33x2_ASAP7_75t_R cut_134 (.A1(req_rdy),
    .A2(\dpath/a_lt_b$in0[6] ),
    .A3(cut_24656),
    .B1(cut_27181),
    .B2(cut_27282),
    .B3(cut_27383),
    .Y(_075_));
 AND2x2_ASAP7_75t_R cut_135 (.A(cut_23343),
    .B(cut_25363),
    .Y(cut_27686));
 OA21x2_ASAP7_75t_R cut_136 (.A1(cut_24454),
    .A2(req_msg[23]),
    .B(cut_24555),
    .Y(cut_27787));
 OA21x2_ASAP7_75t_R cut_137 (.A1(_051_),
    .A2(cut_26777),
    .B(_020_),
    .Y(cut_27484));
 OA21x2_ASAP7_75t_R cut_138 (.A1(_019_),
    .A2(cut_27484),
    .B(_018_),
    .Y(cut_27585));
 XOR2x2_ASAP7_75t_R cut_139 (.A(_050_),
    .B(cut_27585),
    .Y(resp_msg[7]));
 AND3x1_ASAP7_75t_R cut_140 (.A(cut_21222),
    .B(cut_25464),
    .C(resp_msg[7]),
    .Y(cut_27888));
 OA33x2_ASAP7_75t_R cut_141 (.A1(cut_22333),
    .A2(\dpath/a_lt_b$in0[7] ),
    .A3(cut_24656),
    .B1(cut_27686),
    .B2(cut_27787),
    .B3(cut_27888),
    .Y(_076_));
 AND2x2_ASAP7_75t_R cut_142 (.A(cut_23444),
    .B(cut_25363),
    .Y(cut_27989));
 OA21x2_ASAP7_75t_R cut_143 (.A1(cut_24454),
    .A2(req_msg[24]),
    .B(cut_24555),
    .Y(cut_28090));
 XOR2x2_ASAP7_75t_R cut_144 (.A(_016_),
    .B(cut_1999),
    .Y(resp_msg[8]));
 AND3x1_ASAP7_75t_R cut_145 (.A(cut_21222),
    .B(cut_25464),
    .C(resp_msg[8]),
    .Y(cut_28191));
 OA33x2_ASAP7_75t_R cut_146 (.A1(cut_22333),
    .A2(\dpath/a_lt_b$in0[8] ),
    .A3(cut_24656),
    .B1(cut_27989),
    .B2(cut_28090),
    .B3(cut_28191),
    .Y(_077_));
 OA21x2_ASAP7_75t_R cut_147 (.A1(_050_),
    .A2(cut_27585),
    .B(_017_),
    .Y(cut_28292));
 OA21x2_ASAP7_75t_R cut_148 (.A1(_016_),
    .A2(cut_28292),
    .B(_015_),
    .Y(cut_28393));
 XOR2x2_ASAP7_75t_R cut_149 (.A(_049_),
    .B(cut_28393),
    .Y(resp_msg[9]));
 AND3x1_ASAP7_75t_R cut_150 (.A(cut_20717),
    .B(cut_22131),
    .C(resp_msg[9]),
    .Y(cut_28494));
 OA21x2_ASAP7_75t_R cut_151 (.A1(cut_24454),
    .A2(req_msg[25]),
    .B(cut_24555),
    .Y(cut_28595));
 AND2x2_ASAP7_75t_R cut_152 (.A(cut_23545),
    .B(cut_23747),
    .Y(cut_28696));
 OA33x2_ASAP7_75t_R cut_153 (.A1(cut_22333),
    .A2(\dpath/a_lt_b$in0[9] ),
    .A3(cut_24656),
    .B1(cut_28494),
    .B2(cut_28595),
    .B3(cut_28696),
    .Y(_078_));
 AND2x2_ASAP7_75t_R cut_154 (.A(cut_23646),
    .B(cut_25363),
    .Y(cut_28797));
 OA21x2_ASAP7_75t_R cut_155 (.A1(cut_1911),
    .A2(req_msg[26]),
    .B(cut_24353),
    .Y(cut_28898));
 XOR2x2_ASAP7_75t_R cut_156 (.A(_013_),
    .B(cut_20111),
    .Y(resp_msg[10]));
 AND3x1_ASAP7_75t_R cut_157 (.A(cut_21222),
    .B(cut_25464),
    .C(resp_msg[10]),
    .Y(cut_28999));
 OA33x2_ASAP7_75t_R cut_158 (.A1(cut_22333),
    .A2(\dpath/a_lt_b$in0[10] ),
    .A3(cut_22030),
    .B1(cut_28797),
    .B2(cut_28898),
    .B3(cut_28999),
    .Y(_079_));
 AND2x2_ASAP7_75t_R cut_159 (.A(cut_23848),
    .B(cut_25363),
    .Y(cut_292102));
 OA21x2_ASAP7_75t_R cut_160 (.A1(cut_1911),
    .A2(req_msg[27]),
    .B(cut_24353),
    .Y(cut_293103));
 OA21x2_ASAP7_75t_R cut_161 (.A1(_049_),
    .A2(cut_28393),
    .B(_014_),
    .Y(cut_290100));
 OA21x2_ASAP7_75t_R cut_162 (.A1(_013_),
    .A2(cut_290100),
    .B(_012_),
    .Y(cut_291101));
 XOR2x2_ASAP7_75t_R cut_163 (.A(_011_),
    .B(cut_291101),
    .Y(resp_msg[11]));
 AND3x1_ASAP7_75t_R cut_164 (.A(cut_21222),
    .B(cut_25464),
    .C(resp_msg[11]),
    .Y(cut_294104));
 OA33x2_ASAP7_75t_R cut_165 (.A1(cut_22333),
    .A2(\dpath/a_lt_b$in0[11] ),
    .A3(cut_22030),
    .B1(cut_292102),
    .B2(cut_293103),
    .B3(cut_294104),
    .Y(_080_));
 AND2x2_ASAP7_75t_R cut_166 (.A(cut_23949),
    .B(cut_25363),
    .Y(cut_295105));
 OA21x2_ASAP7_75t_R cut_167 (.A1(cut_1911),
    .A2(req_msg[28]),
    .B(cut_24353),
    .Y(cut_296106));
 XOR2x2_ASAP7_75t_R cut_168 (.A(_009_),
    .B(cut_20313),
    .Y(resp_msg[12]));
 AND3x1_ASAP7_75t_R cut_169 (.A(cut_21222),
    .B(cut_25464),
    .C(resp_msg[12]),
    .Y(cut_297107));
 OA33x2_ASAP7_75t_R cut_170 (.A1(cut_22333),
    .A2(\dpath/a_lt_b$in0[12] ),
    .A3(cut_22030),
    .B1(cut_295105),
    .B2(cut_296106),
    .B3(cut_297107),
    .Y(_081_));
 AND2x2_ASAP7_75t_R cut_171 (.A(cut_24050),
    .B(cut_25363),
    .Y(cut_300110));
 OA21x2_ASAP7_75t_R cut_172 (.A1(cut_1911),
    .A2(req_msg[29]),
    .B(cut_24353),
    .Y(cut_301111));
 OA21x2_ASAP7_75t_R cut_173 (.A1(_011_),
    .A2(cut_291101),
    .B(_010_),
    .Y(cut_298108));
 OA21x2_ASAP7_75t_R cut_174 (.A1(_009_),
    .A2(cut_298108),
    .B(_008_),
    .Y(cut_299109));
 XOR2x2_ASAP7_75t_R cut_175 (.A(_007_),
    .B(cut_299109),
    .Y(resp_msg[13]));
 AND3x1_ASAP7_75t_R cut_176 (.A(cut_20717),
    .B(cut_25464),
    .C(resp_msg[13]),
    .Y(cut_302112));
 OA33x2_ASAP7_75t_R cut_177 (.A1(cut_22333),
    .A2(\dpath/a_lt_b$in0[13] ),
    .A3(cut_22030),
    .B1(cut_300110),
    .B2(cut_301111),
    .B3(cut_302112),
    .Y(_082_));
 AND2x2_ASAP7_75t_R cut_178 (.A(cut_24151),
    .B(cut_22232),
    .Y(cut_303113));
 OA21x2_ASAP7_75t_R cut_179 (.A1(cut_1911),
    .A2(req_msg[30]),
    .B(cut_24353),
    .Y(cut_304114));
 XOR2x2_ASAP7_75t_R cut_180 (.A(_005_),
    .B(cut_20515),
    .Y(resp_msg[14]));
 AND3x1_ASAP7_75t_R cut_181 (.A(cut_20717),
    .B(cut_22131),
    .C(resp_msg[14]),
    .Y(cut_305115));
 OA33x2_ASAP7_75t_R cut_182 (.A1(cut_22333),
    .A2(\dpath/a_lt_b$in0[14] ),
    .A3(cut_22030),
    .B1(cut_303113),
    .B2(cut_304114),
    .B3(cut_305115),
    .Y(_083_));
 AND2x2_ASAP7_75t_R cut_183 (.A(cut_24252),
    .B(cut_22232),
    .Y(cut_309119));
 OA21x2_ASAP7_75t_R cut_184 (.A1(cut_1911),
    .A2(req_msg[31]),
    .B(cut_24353),
    .Y(cut_310120));
 OR2x2_ASAP7_75t_R cut_185 (.A(_005_),
    .B(_007_),
    .Y(cut_306116));
 OA21x2_ASAP7_75t_R cut_186 (.A1(_005_),
    .A2(_006_),
    .B(_004_),
    .Y(cut_307117));
 OA21x2_ASAP7_75t_R cut_187 (.A1(cut_299109),
    .A2(cut_306116),
    .B(cut_307117),
    .Y(cut_308118));
 XOR2x2_ASAP7_75t_R cut_188 (.A(_048_),
    .B(cut_308118),
    .Y(resp_msg[15]));
 AND3x1_ASAP7_75t_R cut_189 (.A(cut_20717),
    .B(cut_22131),
    .C(resp_msg[15]),
    .Y(cut_311121));
 OA33x2_ASAP7_75t_R cut_190 (.A1(cut_22333),
    .A2(\dpath/a_lt_b$in0[15] ),
    .A3(cut_22030),
    .B1(cut_309119),
    .B2(cut_310120),
    .B3(cut_311121),
    .Y(_084_));
endmodule
